import lc3b_types::*;

module cache
(

);


cache_datapath cache_datapath
(

);

cache_control cache_control
(
	
);

endmodule : cache
