import lc3b_types::*;

module cache_datapath
(
	// inputs and outputs. 

);

// internal signals



// block assignments. 


endmodule : cache_datapath
